* EESchema Netlist Version 1.1 (Spice format) creation date: sön  1 mar 2015 17:33:45

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
E1  Net-_E1-Pad1_ 0 Net-_C2-Pad1_ Net-_E1-Pad4_ 100		
M1  vd /vg 0 0 nch l=0.18u w=10u		
I1  0 vd DC 500u		
V2  Net-_E1-Pad4_ 0 DC 1		
C2  Net-_C2-Pad1_ 0 1		
R2  Net-_C2-Pad1_ vd 10Mega		
R1  /vg Net-_E1-Pad1_ 10Mega		
C1  /vg Net-_C1-Pad2_ 1		
V1  Net-_C1-Pad2_ 0 DC 0 AC 1		

.include ./models/skew_tt.inc
.include ./models/modelcard3.nmos
.include ./models/modelcard3.pmos

.control
set noaskquit
op
ac dec 10 1 1e9
noise v(vd) V1 dec 10 1 100e9 10
setplot ac1
plot abs(v(vd))
setplot noise1
plot sqrt(inoise_spectrum)
plot db(sqrt(inoise_spectrum))
rusage all
.endc

.end
